--Benjamin Towle
--10/2/2023
--tb_control.vhd
--Used to test our control.vhd module

library IEEE;
use IEEE.std_logic_1164.all;library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.textio.all;             -- For basic I/O

entity tb_control is 
end tb_control;

architecture structure of tb_control is 

component control is 
 port(i_opCode   : in std_logic_vector(5 downto 0); --MIPS instruction opcode (6 bits wide)
	i_funCode  : in std_logic_vector(5 downto 0); --MIPS instruction function code (6 bits wide) used for R-Type instructions
	o_RegDst   : out std_logic;
	o_RegWrite : out std_logic;
	o_memToReg : out std_logic;
	o_memWrite : out std_logic;
	o_ALUSrc   : out std_logic;
	o_ALUOp    : out std_logic_vector(3 downto 0);
	o_signed   : out std_logic;
	o_addSub   : out std_logic;
	o_shiftType : out std_logic;
	o_shiftDir  : out std_logic;
	o_bne       : out std_logic;
	o_beq       : out std_logic;
	o_j         : out std_logic;
	o_jr        : out std_logic;
	o_jal       : out std_logic;
	o_jump      : out std_logic;
	o_branch    : out std_logic);
end component;

signal s_opCode     : std_logic_vector(5 downto 0);
signal s_funCode    : std_logic_vector(5 downto 0);
signal s_RegDst     : std_logic;
signal s_RegWrite   : std_logic;
signal s_memToReg   : std_logic;
signal s_memWrite   : std_logic;
signal s_ALUSrc     : std_logic;
signal s_signed     : std_logic;
signal s_ALUOp      : std_logic_vector(3 downto 0);

signal s_addSub     : std_logic;
signal s_shiftType  : std_logic;
signal s_shiftDir   : std_logic;
signal s_bne        : std_logic;
signal s_beq        : std_logic;
signal s_j          : std_logic;
signal s_jal        : std_logic;
signal s_jr         : std_logic;
signal s_branch     : std_logic;
signal s_jump       : std_logic;

begin 
DUT0: control 

port map(i_opCode   => s_opCode,
	 i_funCode  => s_funCode,
	 o_RegDst   => s_RegDst,
	 o_RegWrite => s_RegWrite,
	 o_memToReg => s_memToReg,
	 o_memWrite => s_memWrite,
	 o_ALUSrc   => s_ALUSrc,
	 o_signed   => s_signed,
	 o_ALUOp    => s_ALUOp, 

	 o_addSub   => s_addSub,
	 o_shiftType => s_shiftType,
	 o_shiftDir  => s_shiftDir,
	 o_bne       => s_bne,
	 o_beq       => s_beq,
	 o_j         => s_j,
	 o_jal       => s_jal,
	 o_jr        => s_jr,
	 o_jump      => s_jump,
	 o_branch    => s_branch);


TEST_CASES: process
begin

s_opCode  <= "000000";
s_funCode <= "010000"; 
wait for 50 ns;   --add instruction

s_opCode  <= "001000";
s_funCode <= "000000"; 
wait for 50 ns;   --addi instruction

s_opCode  <= "000000";
s_funCode <= "100001"; 
wait for 50 ns;   --addu instruction

s_opCode  <= "000000";
s_funCode <= "100100"; 
wait for 50 ns;   --and instruction

s_opCode  <= "001100";
s_funCode <= "000000"; 
wait for 50 ns;   --andi instruction

s_opCode  <= "001111";
s_funCode <= "000000"; 
wait for 50 ns;   --lui instruction

s_opCode  <= "100011";
s_funCode <= "000000"; 
wait for 50 ns;   --lw instruction

s_opCode  <= "000000";
s_funCode <= "100111"; 
wait for 50 ns;   --nor instruction

s_opCode  <= "000000";
s_funCode <= "100110"; 
wait for 50 ns;   --xor instruction

s_opCode  <= "001110";
s_funCode <= "000000"; 
wait for 50 ns;   --xori instruction

s_opCode  <= "000000";
s_funCode <= "100101"; 
wait for 50 ns;   --or instruction

s_opCode  <= "001101";
s_funCode <= "000000"; 
wait for 50 ns;   --ori instruction

s_opCode  <= "000000";
s_funCode <= "101010"; 
wait for 50 ns;   --slt instruction

s_opCode  <= "001010";
s_funCode <= "000000"; 
wait for 50 ns;   --slti instruction

s_opCode  <= "000000";
s_funCode <= "000000"; 
wait for 50 ns;   --sll instruction

s_opCode  <= "000000";
s_funCode <= "000010"; 
wait for 50 ns;   --srl instruction

s_opCode  <= "000000";
s_funCode <= "000011"; 
wait for 50 ns;   --sra instruction

s_opCode  <= "101011";
s_funCode <= "000000"; 
wait for 50 ns;   --sw instruction

s_opCode  <= "000000";
s_funCode <= "100010"; 
wait for 50 ns;   --sub instruction

s_opCode  <= "000000";
s_funCode <= "100011"; 
wait for 50 ns;   --subu instruction

s_opCode  <= "000100";
s_funCode <= "000000"; 
wait for 50 ns;   --beq instruction

s_opCode  <= "000101";
s_funCode <= "000000"; 
wait for 50 ns;   --bne instruction

s_opCode  <= "000010";
s_funCode <= "000000"; 
wait for 50 ns;   --j instruction

s_opCode  <= "000011";
s_funCode <= "000000"; 
wait for 50 ns;   --jal instruction

s_opCode  <= "000000";
s_funCode <= "001000"; 
wait for 50 ns;   --jr instruction

end process;
	  


end structure;