--Benjamin Towle
--11/1/2023
--reg_EX_MEM.vhd
--File contains elements of an N bit register with dffg.vhd as a component

library IEEE;
use IEEE.std_logic_1164.all;

entity reg_EX_MEM is 
   port(i_Flush		 : in std_logic;
		i_CLK        : in std_logic;                          -- Clock input
        i_RST        : in std_logic;                          -- Reset input
        i_WE         : in std_logic;                          -- Write enable input

--INPUTS
	--Control signals used by the MEM stage (input)
	i_memWr      : in std_logic;

	--Control signals forwarded to WB stage (input)
	i_memToReg   : in std_logic;
	i_jal        : in std_logic;
	i_regDst     : in std_logic;
	i_halt       : in std_logic;
	i_regWr      : in std_logic;
	i_Overflow   : in std_logic;
	i_pJPC       : in std_logic_vector(31 downto 0);

	--32-bit and 3-bit inputs
	i_PC_Incremented  : in std_logic_vector(31 downto 0);
	i_RSaddr          : in std_logic_vector(4 downto 0); 
	i_RDaddr          : in std_logic_vector(4 downto 0);
	i_RTaddr          : in std_logic_vector(4 downto 0);
	i_wrAddr          : in std_logic_vector(4 downto 0); 
	i_RTdata          : in std_logic_vector(31 downto 0); 
	i_ALUResult       : in std_logic_vector(31 downto 0);

--OUTPUTS
	--Control signals used by the MEM stage (output)
	o_memWr      : out std_logic;

	--Control signals forwarded to WB stage (output)
	o_memToReg   : out std_logic;
	o_jal        : out std_logic;
	o_regDst     : out std_logic;
	o_halt       : out std_logic;
	o_regWr      : out std_logic;
	o_Overflow   : out std_logic;
	o_pJPC       : out std_logic_vector(31 downto 0); 

	--32-bit and 4-bit outputs
	o_PC_Incremented  : out std_logic_vector(31 downto 0);
	o_RSaddr          : out std_logic_vector(4 downto 0); 
	o_RDaddr          : out std_logic_vector(4 downto 0);
	o_RTaddr          : out std_logic_vector(4 downto 0); 
	o_wrAddr          : out std_logic_vector(4 downto 0); 
	o_RTdata          : out std_logic_vector(31 downto 0);  
	o_ALUResult       : out std_logic_vector(31 downto 0));

end reg_EX_MEM;

architecture structure of reg_EX_MEM is

 component dffg is 
  port(i_CLK        : in std_logic;     -- Clock input
       i_RST        : in std_logic;     -- Reset input
       i_WE         : in std_logic;     -- Write enable input
       i_D          : in std_logic;     -- Data value input
       o_Q          : out std_logic);   -- Data value output
 end component;

 component nBitRegister is 
  generic (N: integer := 32);
   port(i_CLK        : in std_logic;                          -- Clock input
        i_RST        : in std_logic;                          -- Reset input
        i_WE         : in std_logic;                          -- Write enable input
        i_D          : in std_logic_vector(N-1 downto 0);     -- Data value input
        o_Q          : out std_logic_vector(N-1 downto 0));   -- Data value output
 end component;
 
component mux2t1_N is  
	generic(N : integer := 32);
	port(i_S          : in std_logic;
		 i_D0         : in std_logic_vector(N-1 downto 0);
		 i_D1         : in std_logic_vector(N-1 downto 0);
		 o_O          : out std_logic_vector(N-1 downto 0));
end component;

component mux2t1 is
	port(
		i_S	: in std_logic;
		i_D0	: in std_logic;
		i_D1	: in std_logic;
		o_O	: out std_logic);
end component;

signal s_memWr      : std_logic;
signal s_memToReg   : std_logic;
signal s_jal        : std_logic;
signal s_regDst     : std_logic;
signal s_halt       : std_logic;
signal s_regWr      : std_logic;
signal s_Overflow   : std_logic;
signal s_pJPC       : std_logic_vector(31 downto 0);
signal s_PC_Incremented  : std_logic_vector(31 downto 0);
signal s_RSaddr          : std_logic_vector(4 downto 0); 
signal s_RDaddr          : std_logic_vector(4 downto 0);
signal s_RTaddr          : std_logic_vector(4 downto 0);
signal s_WrAddr          : std_logic_vector(4 downto 0); 
signal s_RTdata          : std_logic_vector(31 downto 0); 
signal s_ALUResult       : std_logic_vector(31 downto 0);


begin

--INPUTS
--Control signals used by the MEM stage (input)
	G_memWr : dffg 
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_memWr,
		o_Q    => o_memWr);


	MUX_memWr : mux2t1
		port map(i_S          => i_Flush,
			i_D0         => i_memWr,
			i_D1         => '0',
			o_O          => s_memWr);
	     

	--Control signals forwarded to WB stage (input)
	G_memToReg : dffg 
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_memToReg,
		o_Q    => o_memToReg);

	MUX_memToReg : mux2t1
		port map(i_S          => i_Flush,
			i_D0         => i_memToReg,
			i_D1         => '0',
			o_O          => s_memToReg);
	   
	G_jal : dffg 
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_jal,
		o_Q    => o_jal);

	MUX_jal : mux2t1
		port map(i_S          => i_Flush,
			i_D0         => i_jal,
			i_D1         => '0',
			o_O          => s_jal);
	        
	G_regDst : dffg 
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_regDst,
		o_Q    => o_regDst);

	MUX_regDst : mux2t1
		port map(i_S          => i_Flush,
			i_D0         => i_regDst,
			i_D1         => '0',
			o_O          => s_regDst);
	     
	G_halt : dffg 
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_halt,
		o_Q    => o_halt);

	MUX_halt : mux2t1
		port map(i_S          => i_Flush,
			i_D0         => i_halt,
			i_D1         => '0',
			o_O          => s_halt);
	       
	G_regWr : dffg 
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_regWr,
		o_Q    => o_regWr);

	MUX_regWr : mux2t1
		port map(i_S          => i_Flush,
			i_D0         => i_regWr,
			i_D1         => '0',
			o_O          => s_regWr);

	G_OVFL : dffg 
	port map(i_CLK  => i_CLK,
			 i_RST  => i_RST,
			 i_WE   => i_WE,
			 i_D    => s_Overflow,
			 o_Q    => o_Overflow);

	MUX_OVFL : mux2t1
		port map(i_S          => i_Flush,
			i_D0         => i_Overflow,
			i_D1         => '0',
			o_O          => s_Overflow);
		 

	--32-bit and 3-bit inputs
	G_PC_Incremented : nBitRegister
	generic map (N  => 32)
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_PC_Incremented,
		o_Q    => o_PC_Incremented);


	MUX_PC_Incremented: mux2t1_N
		generic map(N => 32)
		port map(i_S          => i_Flush,
			i_D0         => i_PC_Incremented,
			i_D1         => x"00000000",
			o_O          => s_PC_Incremented);

	G_RSaddr   : nBitRegister
	generic map (N  => 5)
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_RSaddr,
		o_Q    => o_RSaddr);

	MUX_RSaddr: mux2t1_N
		generic map(N => 5)
		port map(i_S          => i_Flush,
			i_D0         => i_RSaddr,
			i_D1         => b"00000",
			o_O          => s_RSaddr);

	G_RDaddr         : nBitRegister
	generic map (N  => 5)
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_RDaddr,
		o_Q    => o_RDaddr);

		
	MUX_RDaddr: mux2t1_N
		generic map(N => 5)
		port map(i_S          => i_Flush,
			i_D0         => i_RDaddr,
			i_D1         => b"00000",
			o_O          => s_RDaddr);

	G_RTaddr         : nBitRegister
	generic map (N  => 5)
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_RTaddr,
		o_Q    => o_RTaddr);


	MUX_RTaddr: mux2t1_N
		generic map(N => 5)
		port map(i_S          => i_Flush,
			i_D0         => i_RTaddr,
			i_D1         => b"00000" ,
			o_O          => s_RTaddr);


	G_WrAddr    : nBitRegister
	generic map (N  => 5)
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_WrAddr,
		o_Q    => o_WrAddr);

	MUX_WrAddr: mux2t1_N
		generic map(N => 5)
		port map(i_S          => i_Flush,
			i_D0         => i_WrAddr,
			i_D1         => b"00000" ,
			o_O          => s_WrAddr);

	G_RTdata   : nBitRegister
	generic map (N  => 32)
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_RTdata,
		o_Q    => o_RTdata);

	MUX_RTdata: mux2t1_N
		generic map(N => 32)
		port map(i_S          => i_Flush,
			i_D0         => i_RTdata,
			i_D1         => x"00000000",
			o_O          => s_RTdata);

	G_ALUResult      : nBitRegister
	generic map (N  => 32)
	port map(i_CLK  => i_CLK,
		i_RST  => i_RST,
		i_WE   => i_WE,
		i_D    => s_ALUResult,
		o_Q    => o_ALUResult);

	MUX_ALUResult: mux2t1_N
		generic map(N => 32)
		port map(i_S          => i_Flush,
			i_D0         => i_ALUResult ,
			i_D1         => x"00000000",
			o_O          => s_ALUResult);
		

	G_pJPC : nBitRegister
	generic map (N => 32) 
	port map(i_CLK  => i_CLK,
			 i_RST  => i_RST,
			 i_WE   => i_WE,
			 i_D    => s_pJPC,
			 o_Q    => o_pJPC);

	MUX_pJPC: mux2t1_N
		generic map(N => 32)
		port map(i_S          => i_Flush,
			i_D0         => i_pJPC,
			i_D1         => x"00000000",
			o_O          => s_pJPC);
	

	
	

end structure;