-------------------------------------------------------------------------
-- Benjamin Towle
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------
-- tb_mux2t1_N.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a testbench for the nbit mux 2t1 unit.
--              
-- 9/4/2023
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.textio.all;             -- For basic I/O

entity tb_mux2t1_N is
 generic(N : integer := 16);
end tb_mux2t1_N;

architecture structure of tb_mux2t1_N is

component mux2t1_N is
  port (i_S : in std_logic;
        i_D0 : in std_logic_vector(N-1 downto 0);
        i_D1 : in std_logic_vector(N-1 downto 0);
        o_O : out std_logic_vector(N-1 downto 0));
end component;


signal s_i_S : std_logic;
signal s_i_D0  : std_logic_vector(N-1 downto 0);
signal s_i_D1   : std_logic_vector(N-1 downto 0);
signal s_o_O   : std_logic_vector(N-1 downto 0);

begin
DUT0: mux2t1_N
port map(i_S     => s_i_S,
	 i_D0    => s_i_D0,
	 i_D1    => s_i_D1,
	 o_O     => s_o_O);



TEST_CASE_1: process
begin

 s_i_S <= '1';
 s_i_D0 <= "1001110000000010";
 s_i_D1 <= "1111011010000011";
--Expect the o_O to be the same as s_i_D1
 

wait for 300 ns;
end process;


end structure;