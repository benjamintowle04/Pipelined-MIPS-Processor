--Benjamin Towle
--10/1/2023
--control.vhd
--To be used to send out all control signals via one module
--More control signals will need to be added to this later, we will keep updating this file as we continue

library IEEE;
use IEEE.std_logic_1164.all;


entity control is 
   port(i_opCode   : in std_logic_vector(5 downto 0); --MIPS instruction opcode (6 bits wide)
	i_funCode  : in std_logic_vector(5 downto 0); --MIPS instruction function code (6 bits wide) used for R-Type instructions
	o_RegDst   : out std_logic;
	o_RegWrite : out std_logic;
	o_memToReg : out std_logic;
	o_memWrite : out std_logic;
	o_ALUSrc   : out std_logic;
	o_ALUOp    : out std_logic_vector(3 downto 0);
	o_signed   : out std_logic;
	o_addSub   : out std_logic;
	o_shiftType : out std_logic;
	o_shiftDir  : out std_logic;
	o_bne       : out std_logic;
	o_beq       : out std_logic;
	o_j         : out std_logic;
	o_jr        : out std_logic;
	o_jal       : out std_logic;
	o_branch    : out std_logic;
	o_jump      : out std_logic;
	o_lui       : out std_logic;
	o_halt      : out std_logic;
	o_ctlExt    : out std_logic);
end control;

architecture behavioral of control is 
begin

process(i_opCode, i_funCode)
begin
  if i_opCode = "000000" then --Case for R-Type instruction
	if i_funCode = "100000" then   --add instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0010"; 
	   o_signed   <= '1';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "100001" then  --addu instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0010"; 
	   o_signed   <= '0';
 	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "100100" then --and instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0011"; 
	   o_signed   <= '0';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "100111" then --nor instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0101"; 
	   o_signed   <= '0';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';  
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "100110" then --xor instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0110"; 
	   o_signed   <= '0';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "100101" then --or instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0111"; 
	   o_signed   <= '0';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "101010" then --slt instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "1000"; 
	   o_signed   <= '1';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "000000" then --sll instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "1001"; 
	   o_signed   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '1';
	   o_addSub   <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "000010" then --srl instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "1001"; 
	   o_signed   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_addSub   <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "000011" then --sra instruction
	   o_RegDst    <= '1';
	   o_RegWrite  <= '1';
	   o_memToReg  <= '0';
	   o_memWrite  <= '0';
	   o_ALUSrc    <= '0';
	   o_ALUOp     <= "1001"; 
	   o_signed    <= '0';
	   o_shiftType <= '1';
	   o_shiftDir  <= '0';
	   o_addSub    <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "100010" then --sub instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0010"; 
	   o_signed   <= '1';
	   o_addSub   <= '1';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "100011" then --subu instruction
	   o_RegDst <= '1';
	   o_RegWrite <= '1';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0010"; 
	   o_signed   <= '0';
	   o_addSub   <= '1';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	elsif i_funCode = "001000" then --jr instruction
	   o_RegDst <= '0';
	   o_RegWrite <= '0';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "1011"; 
	   o_signed   <= '0';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j        <= '0';
	   o_jal      <= '0';
	   o_jr       <= '1';
	   o_jump     <= '1';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	else 
	   o_RegDst <= '0';
	   o_RegWrite <= '0';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0000"; 
	   o_signed   <= '0';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j        <= '0';
	   o_jal      <= '0';
	   o_jr       <= '0';
	   o_jump     <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	end if;


  else  --I and J type instructions
 	if i_opCode = "001000" then --addi instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "0010"; 
	    o_signed   <= '1';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '1';
	elsif i_opCode = "001001" then --addiu instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "0010"; 
	    o_signed   <= '0';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '1';
	elsif i_opCode = "001100" then --andi instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "0011"; 
	    o_signed   <= '0';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '0';
	elsif i_opCode = "001111" then --lui instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "1001"; 
	    o_signed   <= '0';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '1';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '1';
	    o_halt      <= '0';
	    o_ctlExt    <= '0';
	elsif  i_opCode = "100011" then --lw instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '1';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "0010"; 
	    o_signed   <= '0';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '1';
	elsif i_opCode = "001110" then --xori instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "0110"; 
	    o_signed   <= '0';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '0';
	elsif i_opCode = "001101" then --ori instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "0111"; 
	    o_signed   <= '0';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '0';
	elsif i_opCode = "001010" then --slti instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "1000"; 
	    o_signed   <= '1';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '1';
	elsif i_opCode = "101011" then --sw instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '0';
	    o_memToReg <= '0';
	    o_memWrite <= '1';
	    o_ALUSrc   <= '1';
	    o_ALUOp    <= "0010"; 
	    o_signed   <= '0';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '1';
	elsif i_opCode = "000100" then --beq instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '0';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '0';
	    o_ALUOp    <= "0000"; 
	    o_signed   <= '0';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '1';
	    o_branch    <= '1';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '0';
	elsif i_opCode = "000101" then --bne instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '0';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '0';
	    o_ALUOp    <= "0000"; 
	    o_signed   <= '0';
	    o_bne      <= '1';
	    o_beq      <= '0';
	    o_branch   <= '1';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_j         <= '0';   
	    o_jr        <= '0';
	    o_jal       <= '0';
	    o_jump      <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '0';
	elsif i_opCode = "000010" then --j instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '0';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '0';
	    o_ALUOp    <= "1011"; 
	    o_signed   <= '0';
	    o_j        <= '1';
	    o_jal      <= '0';
	    o_jr       <= '0';
	    o_jump     <= '1';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '0';
	elsif i_opCode = "000011" then --jal instruction
	    o_RegDst <= '0';
	    o_RegWrite <= '1';
	    o_memToReg <= '0';
	    o_memWrite <= '0';
	    o_ALUSrc   <= '0';
	    o_ALUOp    <= "1011"; 
	    o_signed   <= '0';
	    o_j        <= '0';
	    o_jal      <= '1';
	    o_jr       <= '0';
	    o_jump     <= '1';
	    o_addSub   <= '0';
	    o_shiftType <= '0';
	    o_shiftDir  <= '0';
	    o_bne       <= '0';
	    o_beq       <= '0';
	    o_branch    <= '0';
	    o_lui       <= '0';
	    o_halt      <= '0';
	    o_ctlExt    <= '0';
	elsif i_opCode = "010100" then --halt instruction 
	   o_RegDst <= '0';
	   o_RegWrite <= '0';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0000"; 
	   o_signed   <= '0';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '1';
	   o_ctlExt    <= '0';
	else 
	   o_RegDst <= '0';
	   o_RegWrite <= '0';
	   o_memToReg <= '0';
	   o_memWrite <= '0';
	   o_ALUSrc   <= '0';
	   o_ALUOp    <= "0000"; 
	   o_signed   <= '0';
	   o_addSub   <= '0';
	   o_shiftType <= '0';
	   o_shiftDir  <= '0';
	   o_bne       <= '0';
	   o_beq       <= '0';
	   o_branch    <= '0';
	   o_j         <= '0';   
	   o_jr        <= '0';
	   o_jal       <= '0';
	   o_jump      <= '0';
	   o_lui       <= '0';
	   o_halt      <= '0';
	   o_ctlExt    <= '0';
	end if;
end if;

end process;





end behavioral;
