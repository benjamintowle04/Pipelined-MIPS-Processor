--Benjamin Towle
--9/11/2023
--tb_nBitDecoder.vhd
--File contains the test bench for my 5 to 32 bit decoder

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.textio.all;  

entity tb_nBitDecoder is 
 generic (N: integer := 5);
end tb_nBitDecoder;

architecture structure of tb_nBitDecoder is 

  component nBitDecoder is 
   port(i_A  : in std_logic_vector(N-1 downto 0);
	o_Q  : out std_logic_vector((2**N) - 1 downto 0));
  end component;

  signal s_i_A  : std_logic_vector(N-1 downto 0);
  signal s_o_Q  : std_logic_vector((2**N) - 1 downto 0); 

begin 
DUT0: nBitDecoder
port map(i_A     => s_i_A,
	 o_Q    => s_o_Q);

 P_TB: process
  begin

s_i_A <= "11111"; --Expect the most significant output bit to be '1'
wait for 100 ns;

s_i_A <= "11010"; --Expect output to be 000001000000000000... (26th bit is set to 1)
wait for 100 ns;

s_i_A <= "00000"; --Expect the least significant bit to be set to 1
wait for 100 ns;
end process;

end structure;