-------------------------------------------------------------------------
-- Benjamin Towle
-- Iowa State University
-------------------------------------------------------------------------
-- tb_nBitRegFile.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a testbench for the Register File
--              
-- 9/15/2023
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.textio.all;             -- For basic I/O

entity tb_nBitRegFile is
generic (
    N : integer := 5;
    gCLK_HPER : time := 50 ns);
end tb_nBitRegFile;

architecture behavior of tb_nBitRegFile is 
-- Calculate the clock period as twice the half-period
constant cCLK_PER  : time := gCLK_HPER * 2;

component nBitRegFile is
   port(i_WA     : in std_logic_vector(N-1 downto 0);
	i_CLK    : in std_logic;
	i_RST    : in std_logic;
	i_DATA   : in std_logic_vector((2**N) - 1 downto 0);
	i_WEN    : in std_logic;
	i_RA1    : in std_logic_vector(N-1 downto 0);
	i_RA2    : in std_logic_vector(N-1 downto 0);
	o_1      : out std_logic_vector((2**N) - 1 downto 0);
	o_2      : out std_logic_vector((2**N) - 1 downto 0));   -- Data value output
end component; 


signal s_WA     :  std_logic_vector(N-1 downto 0);
signal s_CLK    :  std_logic;
signal s_RST    :  std_logic;
signal s_DATA   :  std_logic_vector((2**N) - 1 downto 0);
signal s_WEN    :  std_logic;
signal s_RA1    :  std_logic_vector(N-1 downto 0);
signal s_RA2    :  std_logic_vector(N-1 downto 0);
signal s_o_1    :  std_logic_vector((2**N) - 1 downto 0);
signal s_o_2    :  std_logic_vector((2**N) - 1 downto 0);

begin
DUT0: nBitRegFile

port map (i_WA   => s_WA,
	  i_CLK  => s_CLK,
	  i_RST  => s_RST,
	  i_DATA => s_DATA,
	  i_WEN  => s_WEN,
	  i_RA1  => s_RA1,
	  i_RA2  => s_RA2,
	  o_1    => s_o_1,
	  o_2    => s_o_2);

  --This first process is to setup the clock for the test bench
  --Cycle starts low then goes high
  P_CLK: process
  begin
    s_CLK <= '0';        
    wait for gCLK_HPER; 
    s_CLK <= '1';        
    wait for gCLK_HPER; 
  end process;

TEST_CASES: process
begin

 -- Reset the registers
s_WA   <=  "00000";
s_RST  <=  '1';
s_WEN  <=  '0';
s_DATA <=   x"00000000";
s_RA1  <=   "00000";
s_RA2  <=   "00000";
wait for cCLK_PER;

--Test case 1: store a value in register 0 and read that value in both mux's (o1 and o2)
s_WA    <= "00000";
s_RST   <= '0';
s_WEN   <= '1';
s_DATA  <= x"FEDCBA98";
s_RA1   <= "00000";
s_RA2   <= "00000";
wait for cCLK_PER;


--Test case 2: write a value to register 4 and read that value in o1, then write a value to register 6 and read that value in o2
s_WA    <= "00100";
s_RST   <= '0';
s_WEN   <= '1';
s_DATA  <= x"44444444";
s_RA1   <= "00100";
wait for cCLK_PER;

s_WA    <= "00110";
s_RST   <= '0';
s_WEN   <= '1';
s_DATA  <= x"66666666";
s_RA2   <= "00110";
wait for cCLK_PER;

end process;


end behavior;