-------------------------------------------------------------------------
-- Benjamin Towle
-- Iowa State University
-------------------------------------------------------------------------
-- tb_nBitAdder.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a testbench for the nBitAdder unit.
--              
-- 9/6/2023
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.textio.all;             -- For basic I/O

entity tb_nBitAdder is
 generic(N : integer := 32);
end tb_nBitAdder;

architecture structure of tb_nBitAdder is 
component nBitAdder is
 port(in_A, in_B  : in std_logic_vector(N-1 downto 0);
      in_C        : in std_logic;
      out_S       : out std_logic_vector(N-1 downto 0);
      out_C       : out std_logic);
end component;


signal s_A : std_logic_vector(N-1 downto 0);
signal s_B  : std_logic_vector(N-1 downto 0);
signal s_Cin   : std_logic;
signal s_S   : std_logic_vector(N-1 downto 0);
signal s_Cout   : std_logic;

begin
DUT0: nBitAdder
port map(in_A    => s_A,
	 in_B    => s_B,
	 in_C    => s_Cin,
	 out_S   => s_S,
	 out_C   => s_Cout);



TEST_CASE_1: process
begin

 s_Cin <= '0';
 s_A <= x"";
 s_B <= "";

wait for 300 ns;
end process;


end structure;