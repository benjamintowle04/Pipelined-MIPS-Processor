-------------------------------------------------------------------------
-- Benjamin Towle

-- Iowa State University
-------------------------------------------------------------------------
-- tb_nBitAddSub.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a testbench for the nbit adder/subtracter unit.
--              
-- 9/6/2023
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.textio.all;             -- For basic I/O

entity tb_nBitAddSub is
 generic(N : integer := 32);
end tb_nBitAddSub;

architecture structure of tb_nBitAddSub is 

component nBitAddSub is 
 port(input_A, input_B  : in std_logic_vector(N-1 downto 0);
      nAdd_Sub    : in std_logic;
      output_S    : out std_logic_vector(N-1 downto 0);
      output_C    : out std_logic);
end component;

signal s_input_A, s_input_B  : std_logic_vector(N-1 downto 0);
signal s_nAdd_Sub            : std_logic;
signal s_output_S            : std_logic_vector(N-1 downto 0);
signal s_output_C            : std_logic;


begin
DUT0: nBitAddSub
port map(input_A      => s_input_A,
	 input_B      => s_input_B,
	 nAdd_Sub     => s_nAdd_Sub,
	 output_S     => s_output_S,
	 output_C     => s_output_C);

TEST_CASE_1: process
begin

--$A + $B
 s_input_A     <= x"00080000";
 s_input_B     <= x"00000001"; 
 s_nAdd_Sub <= '1';
wait for 100 ns;

--$A + immediate
 s_input_A     <= x"0000000F";
 s_input_B     <= x"0000000B"; 
 s_nAdd_Sub <= '0';
wait for 100 ns;

--$A - $B
 s_input_A     <= x"0000000F";
 s_input_B     <= x"0000000B"; 
 s_nAdd_Sub <= '1';
wait for 100 ns;

--$A - immediate
 s_input_A     <= x"0000000F";
 s_input_B     <= x"0000000B"; 
 s_nAdd_Sub <= '1';
wait for 100 ns;

end process;


end structure;
